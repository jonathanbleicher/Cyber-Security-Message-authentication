/*------------------------------------------------------------------------------
 * File          : transmitter_manager.sv
 * Project       : RTL
 * Author        : epjoed
 * Creation date : May 24, 2023
 * Description   : 
 *------------------------------------------------------------------------------*/
