/*------------------------------------------------------------------------------
 * File          : receiver_manager.sv
 * Project       : RTL
 * Author        : epjoed
 * Creation date : May 23, 2023
 * Description   : 
 *------------------------------------------------------------------------------*/
